﻿{"Id":null,"Data":{"Id":"e862a319-644a-4b78-a5bb-c3b0fbe4bd52","CounterId":"ed71b345-4af4-44e6-8547-4d10661b6f9a","Timestamp":"2022-09-02T05:37:50.4018654Z","PageSpecificMetrics":null,"Data":182.0},"Metadata":null}