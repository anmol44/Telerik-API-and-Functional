﻿{"Id":null,"Data":{"Id":"19e24df5-0c6e-49e9-ba46-3140f3685c88","CounterId":"7307c8b7-7dd0-414a-8f69-5e44a3031968","Timestamp":"2022-09-02T05:34:44.9857991Z","PageSpecificMetrics":null,"Data":0.0},"Metadata":null}